module imem (input [7:0] Addr , output [15:0] rd);

reg [15:0] RAM[256:0];
initial


begin
RAM[8'b00000000]=16'b0100110000000101;
RAM[8'b00000001]=16'b0100111000001010;
RAM[8'b00000010]=16'b1111110000000000;
RAM[8'b00000011]=16'b1111111000000001;
RAM[8'b00000100]=16'b1011001000000000;
RAM[8'b00000101]=16'b1011010000000001;
RAM[8'b00000110]=16'b0000011011010000;
RAM[8'b00000111]=16'b0100001001111111;
RAM[8'b00001000]=16'b1000001000001010;
RAM[8'b00001001]=16'b0010000000000110;

end



assign rd = RAM[Addr]; 
endmodule